`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/05/2024 02:50:45 PM
// Design Name: 
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 


//////////////////////////////////////////////////////////////////////////////////

module InstMem (input [5:0] addr, output [31:0] data_out);
    reg [31:0] mem [0:63];

    initial begin

//        mem[0] = 32'b000000000000_00000_010_00001_0000011; // lw x1, 0(x0)
//        mem[1] = 32'b000000000100_00000_010_00010_0000011; // lw x2, 4(x0)
//        mem[2] = 32'b000000001000_00000_010_00011_0000011; // lw x3, 8(x0)
        
//              mem[0] = 32'b000000000000_00000_000_00001_0000011; // lb x1, 0(x0)
//              mem[1] = 32'b000000000001_00000_000_00010_0000011; // lb x2, 1(x0)
//              mem[2] = 32'b000000000010_00000_000_00011_0000011; // lb x3, 2(x0)
        
//        mem[3]=32'b0000000_01010_00011_000_00101_0010011; // addi x5, x3, 10     //test addi
//        mem[3] = 32'b0000000_00010_00001_110_00100_0110011; // or x4, x1, x2        
//        mem[4] = 32'b0_000000_00011_00100_000_0100_0_1100011; // beq x4, x3, 4
//        mem[5] = 32'b0000000_00010_00001_000_00011_0110011; // add x3, x1, x2
//        mem[6] = 32'b0000000_00010_00011_000_00101_0110011; // add x5, x3, x2
//        mem[7] = 32'b0000000_00101_00000_010_01100_0100011; // sw x5, 12(x0)
//        mem[8] = 32'b000000001100_00000_010_00110_0000011; // lw x6, 12(x0)
//        mem[9] = 32'b0000000_00001_00110_111_00111_0110011; // and x7, x6, x1
//        mem[10] = 32'b0100000_00010_00001_000_01000_0110011; // sub x8, x1, x2
//        mem[11] = 32'b0000000_00010_00001_000_00000_0110011; // add x0, x1, x2
//        mem[12] = 32'b0000000_00001_00000_000_01001_0110011; // add x9, x0, x1


//////mem[0] = 32'b000000000000_00000_000_00001_0000011; // lb x1, 0(x0)
//////mem[1] = 32'b000000000001_00000_000_00010_0000011; // lb x2, 1(x0)
//mem[2]=32'b00000000001000001000000110110011;   //    add x3, x1, x2       # x3 = x1 + x2
//////mem[2]=32'b00000000100000000000000111101111;// jal x3,8
//////mem[3]=32'b01000000001000001000001000110011;   //    sub x4, x1, x2       # x4 = x1 - x2
//////mem[4]=32'b00000000001000001001001010110011;    //    sll x5, x1, x2       # x5 = x1 << x2
//////mem[5]=32'b00000000001000001101001100110011;     //    srl x6, x1, x2       # x6 = x1 >> x2
//mem[6]=32'b01000000001000001101001110110011;  //    sra x7, x1, x2       # x7 = x1 >> x2 (arithmetic)
//////mem[6]=32'b00000001011000001000011011100111; //jalr x13, 22(x1)
//////mem[7]=32'b00000000001000001111010000110011;   //    and x8, x1, x2       # x8 = x1 & x2
//////mem[8]=32'b00000000001000001110010010110011;   //    or x9, x1, x2        # x9 = x1 | x2
//////mem[9]=32'b00000000001000001100010100110011 ;  //    xor x10, x1, x2      # x10 = x1 ^ x2
//////mem[10]=32'b00000000001000001010010110110011;  //    slt x11, x1, x2      # x11 = (x1 < x2)
//////mem[11]=32'b00000000001000001011011000110011;  //    sltu x12, x1, x2     # x12 = (x1 < x2) (unsigned)

//mem[2] = 32'b00000000101100001000000110010011; // addi x3, x1, 11       # x3 = x1 + 11
//mem[3] = 32'b01000000001000001000001000110011; // subi x4, x1, 11       # x4 = x1 - 11
//mem[4] = 32'b00000000001000001001001010010011; // slli x5, x1, 2        # x5 = x1 << 2
//mem[5] = 32'b00000000001000001101001100010011; // srli x6, x1, 2        # x6 = x1 >> 2
//mem[6] = 32'b01000000001000001101001110010011; // srai x7, x1, 2        # x7 = x1 >> 2 (arithmetic)
//mem[7] = 32'b00000000101100001111010000010011; // andi x8, x1, 11       # x8 = x1 & 11
//mem[8] = 32'b00000000101100001110010010010011; // ori x9, x1, 11        # x9 = x1 | 11
//mem[9] = 32'b00000000101100001100010100010011; // xori x10, x1, 11      # x10 = x1 ^ 11
//mem[10] = 32'b00000000101100001010010110010011; // slti x11, x1, 11      # x11 = (x1 < 11)
//mem[11] = 32'b00000000101100001011011000010011; // sltiu x12, x1, 11     # x12 = (x1 < 11) (unsigned)

//testing lUI and AUIPC
//mem[0] = 32'b00000000000000000010111000110111; //LUI
//mem[1] = 32'b00000000000000000010111000010111; //AUIPC

//testing system calls
mem[0] = 32'b00000000000111111000111110010011; //increment x31
mem[1] = 32'b00000000000111111000111110010011; //increment x31
mem[2] = 32'b00001111111100000000000000001111; //fence
mem[3] = 32'b00000000000111111000111110010011; //increment x31
mem[4] = 32'b00000000000100000000000001110011;//ebreak
mem[5] = 32'b00000000000111111000111110010011; //increment x31
mem[6] = 32'b00000000000000000000000001110011; //ecall
mem[7] = 32'b00000000000111111000111110010011; //increment x31 (should not be executed)




    end

    assign data_out = mem[addr];
endmodule
