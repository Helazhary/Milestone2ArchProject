`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/05/2024 02:50:45 PM
// Design Name: 
// Module Name: InstMem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 


//////////////////////////////////////////////////////////////////////////////////

module InstMem (input [5:0] addr, output [31:0] data_out);
    reg [31:0] mem [0:63];

    initial begin

//        mem[0] = 32'b000000000000_00000_010_00001_0000011; // lw x1, 0(x0)
//        mem[1] = 32'b000000000100_00000_010_00010_0000011; // lw x2, 4(x0)
//        mem[2] = 32'b000000001000_00000_010_00011_0000011; // lw x3, 8(x0)
        
//              mem[0] = 32'b000000000000_00000_000_00001_0000011; // lb x1, 0(x0)
//              mem[1] = 32'b000000000010_00000_001_00010_0000011; // lh x2, 2(x0)
//              mem[2] = 32'b000000000000_00000_010_00011_0000011; // lw x3, 0(x0)
        
      //  mem[3]=32'b0000000_01010_00011_000_00101_0010011; // addi x5, x3, 10     //test addi
//        mem[3] = 32'b0000000_00010_00001_110_00100_0110011; // or x4, x1, x2        
//        mem[4] = 32'b0_000000_00011_00100_000_0100_0_1100011; // beq x4, x3, 4
//        mem[5] = 32'b0000000_00010_00001_000_00011_0110011; // add x3, x1, x2
//        mem[6] = 32'b0000000_00010_00011_000_00101_0110011; // add x5, x3, x2
//        mem[7] = 32'b0000000_00101_00000_010_01100_0100011; // sw x5, 12(x0)
//        mem[8] = 32'b000000001100_00000_010_00110_0000011; // lw x6, 12(x0)
//        mem[9] = 32'b0000000_00001_00110_111_00111_0110011; // and x7, x6, x1
//        mem[10] = 32'b0100000_00010_00001_000_01000_0110011; // sub x8, x1, x2
//        mem[11] = 32'b0000000_00010_00001_000_00000_0110011; // add x0, x1, x2
//        mem[12] = 32'b0000000_00001_00000_000_01001_0110011; // add x9, x0, x1



mem[0] = 32'b00000000000100000000111110010011;
mem[1] = 32'b00000000000000000010000010000011;
mem[2] = 32'b00000000010000000001000100000011;
mem[3] = 32'b00000000100000000000000100000011;
mem[4] = 32'b00000000110000000100001000000011;
mem[5] = 32'b00000001000000000101001010000011;
mem[6] = 32'b00000000001000001000001100110011;
mem[7] = 32'b01000000001000001000001110110011;
mem[8] = 32'b00000000001000001100010000110011;
mem[9] = 32'b00000000001000001110010010110011;
mem[10] = 32'b00000000001000001111010100110011;
mem[11] = 32'b00000000010000001000010110010011;
mem[12] = 32'b00000000010000001100011000010011;
mem[13] = 32'b00000000010000001110011010010011;
mem[14] = 32'b00000000010000001111011100010011;
mem[15] = 32'b00000001111100001101000010110011;
mem[16] = 32'b01000001111100001101000010110011;
mem[17] = 32'b00000000000100001001000010010011;
mem[18] = 32'b00000000000100001101000010010011;
mem[19] = 32'b00000000000000000000001001100011;
mem[20] = 32'b11111111111100001000000010010011;
mem[21] = 32'b00000000000100001000000010010011;
mem[22] = 32'b00000000000100000010000000100011;
mem[23] = 32'b00000000000100000000001000100011;
mem[24] = 32'b00000000000100000001010000100011;


/*
ADDI x31 x0 1 //for incrementing or shifting by 1


LW x1 0(x0)
LH x2 4(x0)
LB x2 8(x0)
LBU x4 12(x0)
LHU x5 16(x0)

ADD x6 x1 x2
SUB x7 x1 x2
XOR x8 x1 x2
OR x9 x1 x2
AND x10 x1 x2


ADDI x11 x1 4
XORI x12 x1 4
ORI x13 x1 4
ANDI x14 x1 4

SRL x1 x1 x31
SRA x1 x1 x31

SLLI x1 x1 1
SRLI x1 x1 1


BEQ x0 x0 4
ADDI x1 x1 -1
ADDI x1 x1 1

SW x1 0(x0)
SB x1 4(x0)
SH x1 8(x0)

*/


    end

    assign data_out = mem[addr];
endmodule
